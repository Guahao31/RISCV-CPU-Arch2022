`ifndef MY_MACROS_VH
`define MY_MACROS_VH

  `define MSTATUS     0
  `define MISA        1
  `define MEDELEG     2
  `define MIDELEG     3
  `define MIE         4
  `define MTVEC       5
  `define MSCRATCH    8
  `define MEPC        9
  `define MCAUSE      10
  `define MTVAL       11

`endif